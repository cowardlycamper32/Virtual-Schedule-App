a,b,1,0
